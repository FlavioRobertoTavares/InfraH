localparam
        RESET   = 0,
        START   = 1,
        ADD     = 2,
        SUB     = 3,
        AND     = 4,
        ANDI    = 5,
        ADDIU   = 6,
        MULT    = 7,
        DIV     = 8,
        JR      = 9,
        MFHI    = 10,
        MFLO    = 11,
        SLL     = 12,
        SLLV    = 13,
        SRA     = 14,
        SRAV    = 15,
        SRL     = 16,
        LUI     = 17,
        SRAM    = 18,
        LB      = 19,
        LH      = 20,
        LW      = 21,
        SB      = 22,
        SH      = 23,
        SW      = 24,
        BNE     = 25,
        BLE     = 26,
        BGT     = 27,
        SLT     = 28,
        SLTI    = 29,
        J       = 30,
        JAL     = 31,
        BREAK   = 31,
        RTE     = 32,
        XCHG    = 33
        ;