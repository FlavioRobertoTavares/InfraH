localparam
        RESET                   = 0 ,
        FETCH                   = 1 ,
        DECODE                  = 2 ,
        OPCODE_INEXISTENTE      = 3 ,
        OVERFLOW                = 4 ,
        DIVZERO                 = 5 ,    
        BREAK                   = 6 ,
        ADD                     = 7 ,
        SUB                     = 8 ,
        AND                     = 9 ,
        ANDI                    = 10,
        ADDIU                   = 11,
        MULT                    = 12,
        DIV                     = 13,
        JR                      = 14,
        MFHI                    = 15,
        MFLO                    = 16,
        SLL                     = 17,
        SLLV                    = 18,
        SRA                     = 19,
        SRAV                    = 20,
        SRL                     = 21,
        LUI                     = 22,
        SRAM                    = 23,
        LB                      = 24,
        LH                      = 25,
        LW                      = 26,
        SB                      = 27,
        SH                      = 28,
        SW                      = 29,
        BNE                     = 30,
        BLE                     = 31,
        BGT                     = 32,
        BEQ                     = 33,
        SLT                     = 34,
        SLTI                    = 35,
        J                       = 36,
        JAL                     = 37,
        RTE                     = 38,
        XCHG                    = 39,
        ADDI                    = 40
        ;