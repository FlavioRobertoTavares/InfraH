integer i = 0;
localparam  
    RESET   = i++,
    START   = i++,
    ADD     = i++,
    SUB     = i++,
    AND     = i++,
    ANDI    = i++,
    ADDIU   = i++,
    MULT    = i++,
    DIV     = i++,
    JR      = i++,
    MFHI    = i++,
    MFLO    = i++,
    SLL     = i++,
    SLLV    = i++,
    SRA     = i++,
    SRAV    = i++,
    SRL     = i++,
    LUI     = i++,
    SRAM    = i++,
    LB      = i++,
    LH      = i++,
    LW      = i++,
    SB      = i++,
    SH      = i++,
    SW      = i++,
    BNE     = i++,
    BLE     = i++,
    BGT     = i++,
    SLT     = i++,
    SLTI    = i++,
    J       = i++,
    JAL     = i++,
    BREAK   = i++,
    RTE     = i++,
    XCHG    = i++
    ;