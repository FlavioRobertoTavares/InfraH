module Controle #(
    
) (
    ports
);
    
endmodule