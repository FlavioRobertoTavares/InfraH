`include "Estados.vh"

module Controle (
    
);
    
endmodule