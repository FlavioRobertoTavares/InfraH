module Controle (
   
);
    `include "Estados.vh"
endmodule