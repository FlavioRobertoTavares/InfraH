localparam
        RESET                   = 0 ,
        FETCH                   = 1 ,
        DECODE                  = 2 ,
        OPCODE_INEXISTENTE      = 3 ,
        OVERFLOW                = 4 ,
        DIVZERO                 = 5 ,    
        BREAK                   = 6 ,
        ADD                     = 7 ,
        SUB                     = 8 ,
        AND                     = 9 ,
        ANDI                    = 10,
        ADDIU                   = 11,
        MULT                    = 12,
        DIV                     = 13,
        JR                      = 14,
        MFHI                    = 15,
        MFLO                    = 16,
        SLL                     = 17,
        SLLV                    = 18,
        SRA                     = 19,
        SRAV                    = 20,
        SRL                     = 21,
        LUI                     = 22,
        SRAM                    = 23,
        MEM                     = 24,
        LB                      = 25,
        LH                      = 26,
        LW                      = 27,
        SB                      = 28,
        SH                      = 29,
        SW                      = 30,
        BNE                     = 31,
        BLE                     = 32,
        BGT                     = 33,
        BEQ                     = 34,
        SLT                     = 35,
        SLTI                    = 36,
        J                       = 37,
        JAL                     = 38,
        RTE                     = 39,
        XCHG                    = 40,
        ADDI                    = 41,
        ADDI_WRITE              = 42
        ;